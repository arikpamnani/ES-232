module decoder(input en, input [3:0] in, output [15:0] out);
	
	reg out;
	always @ (en, in)
	begin
		if(en)	
			begin
				case(in)
					4'b0000 : out = 16'b0000000000000001;
					4'b0001 : out = 16'b0000000000000010;
					4'b0010 : out = 16'b000000000000010;
					4'b0011 : out = 16'b000000000000100;
					4'b0100 : out = 16'b000000000001000;
					4'b0101 : out = 16'b000000000010000;
					4'b0110 : out = 16'b000000000100000;
					4'b0111 : out = 16'b000000001000000;
					4'b1000 : out = 16'b000000010000000;
					4'b1001 : out = 16'b000000100000000;
					4'b1010 : out = 16'b000001000000000;
					4'b1011 : out = 16'b000010000000000;
					4'b1100 : out = 16'b000100000000000;
					4'b1101 : out = 16'b001000000000000;
					4'b1110 : out = 16'b010000000000000;
					4'b1111 : out = 16'b100000000000000;	
				endcase
			end
		else
			out = 16'b0000000000000000;
	end
	
endmodule
